`timescale 1ns/1ps

module alu_test;

reg [31:0] regA,regB;
reg [31:0] instruction;

wire [2:0] flags;
wire [31:0] result;


alu testalu(instruction, regA, regB, result, flags);

initial
begin

$display("     instruction :op :func:   regA   :  regB   : result  :flags");
$monitor("%s   %h :%h : %h : %h :%h :%h :  %b",
testalu.reg_str, instruction, testalu.opcode, testalu.func, regA , regB, result, flags);

// add (overflow)
#10 instruction <= 32'b0000_0000_0010_0000_0001_1000_0010_0000;
regA <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;


// add 
#10 instruction <= 32'b0000_0000_0010_0000_0001_1000_0010_0000;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;

// addu (overflow)
#10 instruction <= 32'b0000_0000_0010_0000_0001_1000_0010_0001;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;


// addu
#10 instruction <= 32'b0000_0000_0010_0000_0001_1000_0010_0001;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1110;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;


// addi (overflow)
#10 instruction <= 32'b0010_0000_0000_0000_0000_0000_0000_0001; //regA = rs
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;


// addi
#10 instruction <= 32'b0010_0000_0010_0000_0000_0000_0000_0001; //regB = rs
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001; 

// addiu (overflow)
#10 instruction <= 32'b0010_0100_0010_0000_1111_1111_1111_1111; 
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001; 

// addiu
#10 instruction <= 32'b0010_0100_0010_0000_1000_0000_0000_0001; 
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001; 

// and
#10 instruction <= 32'b0000_0000_0010_0000_0001_1000_0010_0100;
regA <= 32'b0101_1010_0000_1101_1101_1101_1101_1101;
regB <= 32'b1010_0101_1111_0010_0010_0010_0010_0011;       // result should be 1


// andi
#10 instruction <= 32'b0011_0000_0000_0000_1000_0000_0000_0000;  // imme = 1000_0000_0000_0000 should be -> 0000_0000_0000_0000_1000_0000_0000_0000 
regA <= 32'b1111_1111_1111_1111_1000_0000_1101_1101;
regB <= 32'b1010_0101_1111_0010_0010_0010_0010_0011;      // not used, result should be 0000 8000

// nor
#10 instruction <= 32'b0000_0000_0010_0000_0001_1000_0010_0111;
regA <= 32'b0111_1111_1111_1111_1111_1111_1111_1110;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;      //result should be 1


// or
#10 instruction <= 32'b0000_0000_0010_0000_0001_1000_0010_0101;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
regB <= 32'b1111_1111_1111_1111_1111_1111_1111_0001;     // result should be ffff fff1


// ori
#10 instruction <= 32'b0011_0100_0000_0000_1000_0000_0000_0001;  // imme = 1000_0000_0000_0001 should be -> 0000_0000_0000_0000_1000_0000_0000_0001
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
regB <= 32'b1111_1111_1111_1111_1111_1111_1111_0001;            // result should be 0000 8001

// sll
#10 instruction <= 32'b0000_0000_0000_0000_0001_0010_0000_0000;
regA <= 32'b0000_0000_0000_0000_0000_0001_0000_0000;             // result should be 0001 0000
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001; 

// sllv
#10 instruction<=32'b0000_0000_0000_0001_0001_0000_0000_0100;
regA <= 32'b1111_1101_1101_1101_1101_1101_1100_1000;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;            // result should be 0000 0100


// sra
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_1100_0011;
regA <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;           // result should be f000 0000


// srav
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0000_0111;
regA <= 32'b1101_1101_1101_1101_1101_1101_1100_0111;  
regB <= 32'b1000_0000_0000_0000_0000_0000_0111_1111;          // result should be ff00 0000


// srl
#10 instruction <= 32'b0000_0000_0000_0001_0001_0001_1100_0010;
regA <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;
regB <= 32'b1000_0000_0000_0000_0000_0000_0111_1111;         // result should be 0100 0000


// srlv
#10 instruction<=32'b0000_0000_0000_0001_0001_0000_0000_0110;
regA<=32'b1101_1101_1101_1101_1101_1101_1100_0011;
regB<=32'b1000_0000_0000_0000_0000_0000_0000_0111;           // result should be 1000 0000


// sub
#10 instruction<=32'b0000_0000_0000_0001_0001_1000_0010_0010;
regA<=32'b0110_1101_1101_1101_1101_1101_1101_1101;
regB<=32'b1000_0000_0000_0000_0000_0000_0000_0001;          // should be an overflow


// subu
#10 instruction <= 32'b0000_0000_0010_0000_0001_1000_0010_0011;
regA<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB<=32'b0000_0000_0000_0000_0000_0000_0000_0001;          // result should be 2


// xor
#10 instruction<=32'b0000_0000_0010_0000_0001_1000_0010_0110;
regA<=32'b0110_1101_1101_1101_1101_1101_1101_1101;
regB<=32'b1001_0010_0010_0010_0010_0010_0010_0010;          // result should be ffff ffff             


// xori
#10 instruction<=32'b0011_1000_0000_0001_1000_0000_0000_1111;   // imme -> 0000 0000 0000 0000 1000 0000 0000 1111
regA<=32'b0000_0000_0000_0000_1000_0000_0000_0000;              // result should be 0000 000f


// slt
#10 instruction<=32'b0000_0000_0010_0000_0001_1000_0010_1010;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;            // negative flag


// sltu
#10 instruction<=32'b0000_0000_0010_0000_0001_1000_0010_1011;
regA<=32'b1110_1101_1101_1101_1101_1101_1101_1101;
regB<=32'b0000_0000_0000_0000_0000_0000_0000_0001;             // negative flag  


// slti
#10 instruction<=32'b0010_1000_0010_0000_0001_1000_0010_1011;
regA<=32'b0110_1101_1101_1101_1101_1101_1101_1101;
regB<=32'b1000_0000_0000_0000_0000_0000_0000_0001;            // negative flag


// sltiu
#10 instruction<=32'b0010_1100_0010_0000_1001_1000_0010_1011;
regA<=32'b0110_1101_1101_1101_1101_1101_1101_1101;
regB<=32'b1000_0000_0000_0000_0000_0000_0000_0001;            // negative flag

// beq
#10 instruction<=32'b0001_0000_0010_0000_0001_1000_0010_1011;
regA<=32'b0110_1101_1101_1101_1101_1101_1101_1101;
regB<=32'b0110_1101_1101_1101_1101_1101_1101_1101;                     // zero flag

// beq
#10 instruction<=32'b0001_0000_0010_0000_0001_1000_0010_1011;
regA<=32'b0110_1101_1101_1101_1101_1101_1101_1101;
regB<=32'b0110_1101_1101_1101_1101_1101_1101_1100;                     // no flag

// bne
#10 instruction<=32'b0001_0100_0010_0000_0001_1000_0010_1011;
regA<=32'b0110_1101_1101_1101_1101_1101_1101_1101;
regB<=32'b0110_1101_1101_1101_1101_1101_1101_1101;                    // zero flag

// bne
#10 instruction<=32'b0001_0100_0010_0000_0001_1000_0010_1011;
regA<=32'b0110_1101_1101_1101_1101_1101_1101_1101;
regB<=32'b0110_1101_1101_1101_1101_1101_1101_1100;                    // no flag

// lw
#10 instruction <= 32'b1000_1100_0000_0001_1001_1001_1001_1000;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_1111;                 // result should be ffff9999

// sw
#10 instruction <= 32'b1010_1100_0000_0001_1001_1001_1001_1000;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_1111;                 // result should be ffff9999

#10 $finish;
end
endmodule